`include "src/sysarr.v"

module tb_sysarr();

reg [31:0] l11, l21, l31, l41, u11, u12, u13, u14;
wire [31:0] r11, r12, r13, r14, r21, r22, r23, r24, r31, r32, r33, r34, r41, r42, r43, r44;

sysarr uut(
    l11, l21, l31, l41, u11, u12, u13, u14,
    clk, rst,
    r11, r12, r13, r14, r21, r22, r23, r24, r31, r32, r33, r34, r41, r42, r43, r44
);

reg rst = 1'b0;
reg clk = 1'b1;
always #5 clk = ~clk;

initial begin
    rst <= 1'b1;

    @(posedge clk);

    rst <= 1'b0;

    //A -> identity, B -> identity, C -> identity
    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    wait_sysarr();
    stat();
    rst <= 1'b1;

    @(posedge clk);

    rst <= 1'b0;

    //A -> 1, B -> 1, C -> 4
    l11 <= 32'h3f800000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h3f800000;

    wait_sysarr();
    stat();

    $finish;
end

task wait_sysarr(); begin
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
end
endtask
task stat(); begin
    $display("");
    $display("%h %h %h %h\n%h %h %h %h\n%h %h %h %h\n%h %h %h %h",
        r11, r12, r13, r14,
        r21, r22, r23, r24,
        r31, r32, r33, r34,
        r41, r42, r43, r44
    );
end
endtask
endmodule
