`include "src/sysarr.v"

module tb_sysarr();

reg [31:0] l11, l21, l31, l41, u11, u12, u13, u14;
wire [4:0] count;

sysarr uut(l11, l21, l31, l41, u11, u12, u13, u14,
    clk, rst, count);

reg rst = 1'b0;
reg clk = 1'b1;
always #5 clk = ~clk;

initial begin
    rst <= 1'b1;

    @(posedge clk);

    rst <= 1'b0;

    //A -> identity, B -> identity, C -> identity
    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    wait_sysarr();
    stat();
    rst <= 1'b1;

    @(posedge clk);

    rst <= 1'b0;

    //A -> 1, B -> 1, C -> 4
    l11 <= 32'h3f800000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h00000000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h00000000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h00000000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h00000000;

    @(posedge clk);

    l11 <= 32'h3f800000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h3f800000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h3f800000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h3f800000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h3f800000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h3f800000;
    u14 <= 32'h3f800000;

    @(posedge clk);

    l11 <= 32'h00000000;
    l21 <= 32'h00000000;
    l31 <= 32'h00000000;
    l41 <= 32'h3f800000;

    u11 <= 32'h00000000;
    u12 <= 32'h00000000;
    u13 <= 32'h00000000;
    u14 <= 32'h3f800000;

    wait_sysarr();
    stat();

    $finish;
end

task wait_sysarr(); begin
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
    @(posedge clk);
end
endtask
task stat(); begin
    $display("");
    $display("count: %d\n%h %h %h %h\n%h %h %h %h\n%h %h %h %h\n%h %h %h %h",
        uut.count,
        uut.r11, uut.r12, uut.r13, uut.r14,
        uut.r21, uut.r22, uut.r23, uut.r24,
        uut.r31, uut.r32, uut.r33, uut.r34,
        uut.r41, uut.r42, uut.r43, uut.r44
    );
end
endtask
endmodule
